library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity asd is

end;

architecture asdf of asd is
begin

end asdf;

